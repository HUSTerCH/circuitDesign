** Profile: "SCHEMATIC1-MOSFET_TRAN"  [ D:\Desktop\StudyAndWork\circuitDesgin\CircuitDesignExperiment_lc\2\MOSFET-PSpiceFiles\SCHEMATIC1\MOSFET_TRAN.sim ] 

** Creating circuit file "MOSFET_TRAN.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/OrCAD/OrCAD_16.6_Lite/tools/pspice/library/pwrmos.lib" 
* From [PSPICE NETLIST] section of D:\SPB_data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 4ms 0 1us 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
